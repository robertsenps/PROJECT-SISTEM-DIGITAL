LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY bcd IS PORT (
  SW    : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
  HEX1  : OUT STD_LOGIC_VECTOR (1 TO 7);
  HEX2	: OUT STD_LOGIC_VECTOR (1 TO 7));
END bcd;

ARCHITECTURE behavioral OF bcd IS

  CONSTANT NOL      : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
  CONSTANT SATU     : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
  CONSTANT DUA      : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
  CONSTANT TIGA     : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
  CONSTANT EMPAT    : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
  CONSTANT LIMA     : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
  CONSTANT ENAM     : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
  CONSTANT TUJUH    : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";
  CONSTANT DELAPAN  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
  CONSTANT SEMBILAN : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
  CONSTANT SEPULUH	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";

BEGIN
  
  PROCESS(SW)
  BEGIN
  CASE SW IS    -- Active LOW
  WHEN NOL      => HEX1 <= "0000001"; HEX2 <= "0000001";
  WHEN SATU     => HEX1 <= "1001111"; HEX2 <= "0000001";
  WHEN DUA      => HEX1 <= "0010010"; HEX2 <= "0000001";
  WHEN TIGA     => HEX1 <= "0000110"; HEX2 <= "0000001";
  WHEN EMPAT    => HEX1 <= "1001100"; HEX2 <= "0000001";
  WHEN LIMA     => HEX1 <= "0100100"; HEX2 <= "0000001";
  WHEN ENAM     => HEX1 <= "0100000"; HEX2 <= "0000001";
  WHEN TUJUH    => HEX1 <= "0001111"; HEX2 <= "0000001";
  WHEN DELAPAN  => HEX1 <= "0000000"; HEX2 <= "0000001";
  WHEN SEMBILAN => HEX1 <= "0000100"; HEX2 <= "0000001";
  WHEN SEPULUH	=> HEX1 <= "0000001"; HEX2 <= "1001111";
  WHEN OTHERS   => HEX1 <= "1111111"; HEX2 <= "1111111";
  END CASE;
  END PROCESS;

END behavioral;